library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package configpkg is
	constant rows: integer := 0;
	constant columns: integer := 1;
	constant size_opcode: integer := 0;
	constant size_address: integer := 0;
	constant size_instr: integer := 0;


	constant size_UROM: integer := 0;
	constant size_UROM_address: integer := 0;
	constant size_UROM_instruction: integer := 0;
	constant number_of_urom_instructions: integer := 0;


end configpkg;
